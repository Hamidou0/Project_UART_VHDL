library verilog;
use verilog.vl_types.all;
entity right8_vlg_vec_tst is
end right8_vlg_vec_tst;
