library verilog;
use verilog.vl_types.all;
entity upcounter_8b_vlg_vec_tst is
end upcounter_8b_vlg_vec_tst;
