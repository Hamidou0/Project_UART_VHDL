library verilog;
use verilog.vl_types.all;
entity baude_gen_vlg_vec_tst is
end baude_gen_vlg_vec_tst;
