library verilog;
use verilog.vl_types.all;
entity left8_vlg_vec_tst is
end left8_vlg_vec_tst;
