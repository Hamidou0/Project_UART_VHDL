library verilog;
use verilog.vl_types.all;
entity baude_gen_vlg_check_tst is
    port(
        clock_41        : in     vl_logic;
        clock_Hz        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end baude_gen_vlg_check_tst;
